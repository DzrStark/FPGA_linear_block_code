library verilog;
use verilog.vl_types.all;
entity hanming_decode_mif_vlg_tst is
end hanming_decode_mif_vlg_tst;
