library verilog;
use verilog.vl_types.all;
entity divider7 is
    port(
        clk             : in     vl_logic;
        clk_out         : out    vl_logic
    );
end divider7;
